-- i2c_si53304.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity i2c_si53304 is
	port (
		bladerf_oc_i2c_master_0_clock_sink_clk           : in  std_logic := '0'; --  bladerf_oc_i2c_master_0_clock_sink.clk
		bladerf_oc_i2c_master_0_conduit_end_scl_pad_o    : out std_logic;        -- bladerf_oc_i2c_master_0_conduit_end.scl_pad_o
		bladerf_oc_i2c_master_0_conduit_end_scl_padoen_o : out std_logic;        --                                    .scl_padoen_o
		bladerf_oc_i2c_master_0_conduit_end_sda_pad_i    : in  std_logic := '0'; --                                    .sda_pad_i
		bladerf_oc_i2c_master_0_conduit_end_sda_pad_o    : out std_logic;        --                                    .sda_pad_o
		bladerf_oc_i2c_master_0_conduit_end_sda_padoen_o : out std_logic;        --                                    .sda_padoen_o
		bladerf_oc_i2c_master_0_conduit_end_arst_i       : in  std_logic := '0'; --                                    .arst_i
		bladerf_oc_i2c_master_0_conduit_end_scl_pad_i    : in  std_logic := '0'; --                                    .scl_pad_i
		bladerf_oc_i2c_master_0_reset_sink_reset         : in  std_logic := '0'  --  bladerf_oc_i2c_master_0_reset_sink.reset
	);
end entity i2c_si53304;

architecture rtl of i2c_si53304 is
	component i2c_master_top is
		generic (
			ARST_LVL : integer := 0
		);
		port (
			wb_clk_i     : in  std_logic                    := 'X';             -- clk
			wb_rst_i     : in  std_logic                    := 'X';             -- reset
			scl_pad_o    : out std_logic;                                       -- scl_pad_o
			scl_padoen_o : out std_logic;                                       -- scl_padoen_o
			sda_pad_i    : in  std_logic                    := 'X';             -- sda_pad_i
			sda_pad_o    : out std_logic;                                       -- sda_pad_o
			sda_padoen_o : out std_logic;                                       -- sda_padoen_o
			arst_i       : in  std_logic                    := 'X';             -- arst_i
			scl_pad_i    : in  std_logic                    := 'X';             -- scl_pad_i
			wb_inta_o    : out std_logic;                                       -- irq
			wb_dat_i     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o     : out std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i      : in  std_logic                    := 'X';             -- write
			wb_stb_i     : in  std_logic                    := 'X';             -- byteenable
			wb_cyc_i     : in  std_logic                    := 'X';             -- chipselect
			wb_ack_o     : out std_logic;                                       -- waitrequest_n
			wb_adr_i     : in  std_logic_vector(2 downto 0) := (others => 'X')  -- address
		);
	end component i2c_master_top;

begin

	bladerf_oc_i2c_master_0 : component i2c_master_top
		generic map (
			ARST_LVL => 1
		)
		port map (
			wb_clk_i     => bladerf_oc_i2c_master_0_clock_sink_clk,           --            clock_sink.clk
			wb_rst_i     => bladerf_oc_i2c_master_0_reset_sink_reset,         --            reset_sink.reset
			scl_pad_o    => bladerf_oc_i2c_master_0_conduit_end_scl_pad_o,    --           conduit_end.scl_pad_o
			scl_padoen_o => bladerf_oc_i2c_master_0_conduit_end_scl_padoen_o, --                      .scl_padoen_o
			sda_pad_i    => bladerf_oc_i2c_master_0_conduit_end_sda_pad_i,    --                      .sda_pad_i
			sda_pad_o    => bladerf_oc_i2c_master_0_conduit_end_sda_pad_o,    --                      .sda_pad_o
			sda_padoen_o => bladerf_oc_i2c_master_0_conduit_end_sda_padoen_o, --                      .sda_padoen_o
			arst_i       => bladerf_oc_i2c_master_0_conduit_end_arst_i,       --                      .arst_i
			scl_pad_i    => bladerf_oc_i2c_master_0_conduit_end_scl_pad_i,    --                      .scl_pad_i
			wb_inta_o    => open,                                             --      interrupt_sender.irq
			wb_dat_i     => open,                                             -- bladerf_oc_i2c_master.writedata
			wb_dat_o     => open,                                             --                      .readdata
			wb_we_i      => open,                                             --                      .write
			wb_stb_i     => open,                                             --                      .byteenable
			wb_cyc_i     => open,                                             --                      .chipselect
			wb_ack_o     => open,                                             --                      .waitrequest_n
			wb_adr_i     => open                                              --                      .address
		);

end architecture rtl; -- of i2c_si53304
